
module cordic (
    input clk,
    input rst_n,
    input start,
    input [15:0] angle,
    output reg [15:0] cos,
    output reg [15:0] sin
);

endmodule